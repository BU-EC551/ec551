`timescale 1ns / 1ps
module orgate(a,b,c
    );
	input a;
	input b;
	output c;
	or o1(c,a,b);

endmodule
